package rr is
	constant N:natural:=1;
end rr;

