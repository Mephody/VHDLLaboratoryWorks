package types is
	type mili_in_type is (z1, z2, z3);
	type mili_out_type is (w1, w2, w3, w4, w5);
	type T_state is (a1, a2, a3, a4);
end;
