package pack is
	constant n:natural:=10;
	type ai is array (1 to n) of integer;
end;
